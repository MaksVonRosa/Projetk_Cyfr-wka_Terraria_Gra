module draw_char (
    input  logic clk,
    input  logic rst,
    input  logic stepleft,
    input  logic stepright,
    input  logic stepjump,
    input  logic on_ground,
    input  logic mouse_left,
    output logic [11:0] pos_x_out, pos_y_out,


    vga_if.in  vga_char_in,
    vga_if.out vga_char_out,

    vga_if.in  vga_wpn_in
    //vga_if.out  vga_wpn_out

    
);

    // logic [11:0] pos_x, pos_y;
    assign pos_x_out = pos_x;
    assign pos_y_out = pos_y;
    logic flip_h;

    logic draw_weapon;

    // Character Movement
    char_ctrl u_ctrl (
        .clk(clk),
        .rst(rst),
        .stepleft(stepleft),
        .stepright(stepright),
        .stepjump(stepjump),
        .on_ground(on_ground),
        .pos_x(pos_x),
        .pos_y(pos_y),
        .flip_h(flip_h),
        .draw_weapon(draw_weapon),
        .mouse_left(mouse_left)
    );

    // Character Draw
    char_draw u_draw (
        .clk(clk),
        .rst(rst),
        .pos_x(pos_x),
        .pos_y(pos_y),
        .flip_h(flip_h),
        .vga_in(vga_char_in),
        .vga_out(vga_wpn_in)
    );
    wpn_draw_def u_wpn_draw_def (
        .clk(clk),
        .rst(rst),
        .pos_x(pos_x),
        .pos_y(pos_y),
        .draw_enable(draw_weapon),
        .flip_h(flip_h),
        .vga_in(vga_wpn_in),
        .vga_out(vga_char_out)
    );

endmodule
